module top_module
(
    
    input [39:0] a1,b1,
    output [77:0] c1
   
);
  assign c1 = a1*b1;

endmodule
