module top_module
(
    
    input a1,b1,
    output [1:0] c1
   
);
  assign c1 = a1*b1;


endmodule
